// Code your design here
///////////////////////////////////////////////////////////////////////////

//
// File name   : mux.sv
// Title       : MUX module 
// Project     : SystemVerilog Training

// Description : Defines the mux module 
// Notes       :
//
///////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ns

module mux
(
  input  logic       clock  ,
  input  logic [3:0] ip1    ,
  input  logic [3:0] ip2    ,
  input  logic [3:0] ip3    ,
  input  logic       sel1   ,
  input  logic       sel2   ,
  input  logic       sel3   ,
  output logic [3:0] mux_op  
) ;

always @(posedge clock)
  if (sel1 == 1)
    mux_op <= ip1 ;
  else
    if (sel2 == 1)
      mux_op <= ip2 ;
    else
      if (sel3 == 1)
        mux_op <= ip3 ;
  
    
// assertions go here
//#### edit ###
  
   //----------------------//
  
  property P1;
    @(posedge clock)
    sel1 |=> (mux_op == $past(ip1, 1));
    endproperty
  
  
  property P2;
    @(posedge clock)
    ((sel1 == 1'b0) & (sel2 == 1'b1)) |=> (mux_op == $past(ip2, 1));
    endproperty
  
  
  property P3;
    @(posedge clock)
    ((sel1 == 1'b0) & (sel2 == 1'b0) & (sel3 == 1'b1)) |=> (mux_op == $past(ip3, 1));
    endproperty
  
  
  SEL1_assertion : assert property (P1)
    $display ("###------Congrats!------### SEL1_asseration passed ### : %0t", $time);
    else $fatal("###----------Attentation SEL1_asseration Failed--------### : %0t", $time);
  
    
    
   
    SEL2_assertion : assert property (P2)
      $display ("###------Congrats!------### SEL2_asseration passed ### : %0t", $time);
      else $fatal("###----------Attentation SEL2_asseration Failed--------### : %0t", $time);
  
  
      
      
      SEL3_assertion : assert property (P3)
        $display ("###------Congrats!------### SEL3_asseration passed ### : %0t", $time);
        else $fatal("###----------Attentation SEL3_asseration Failed--------### : %0t", $time);
  
    
    
    //-------------------//



//#### end of edit ###
endmodule
