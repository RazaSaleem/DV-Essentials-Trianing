// Code your design here
module register # (parameter WIDTH=8) (data_in, load, clk, rst, data_out);
  input	wire clk  ;
  input wire rst  ;
  input wire load ;
  input wire [WIDTH-1:0] data_in;
  output reg [WIDTH-1:0] data_out;
  
  always @(posedge clk)
    if( rst )
      data_out <= 0;
  else if (load)
    data_out <=data_in;
  else
    data_out <= data_out;
 endmodule
